module shift(
	input logic [7:0] A, B,
	input logic [7:0] X,
	output logic [7:0] new_A, new_B
);



endmodule 