module adder_9(
	input logic [8:0] XA, S, //S is sign-extended switches
	output logic [7:0] OUT
);



endmodule 